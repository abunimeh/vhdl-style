-- This file is encoded
-- using DOS convention
-- That is \r\n
